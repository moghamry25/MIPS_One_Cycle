module Control_Unit(
    port_list
);
    
endmodule